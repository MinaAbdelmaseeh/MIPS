-----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/01/2022 08:15:00 PM
-- Design Name: 
-- Module Name: MIPS_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MIPS_tb is
--  Port ( );
end MIPS_tb;


architecture Behavioral of MIPS_tb is
component MIPS
port(
    clk: in STD_LOGIC
    );
end component;

signal clk : std_logic;
begin
processor: MIPS port map(clk);

process
begin
clk<='0';   wait for 10 ns;
clk<='1';   wait for 10 ns;
end process;

end Behavioral;
